`default_nettype none
`include "primitives.v"
`include "data_phy.v"
`include "clock_alignment.v"
`include "output_clock.v"


module syzygy_adc #(
    parameter ARCHITECTURE = "7-series",
    parameter OUTPUT_CLOCK = 1,
    parameter IOSTANDARD = "LVDS_25",
    parameter BUFR_DIVIDE_CLOCK = "4"
) (
    input wire clk,
    input wire idelay_ref,  //200mhz
    input wire async_rst,

    //ADC physical pins
    input wire [1:0] adc0_p, adc0_n,    
    input wire [1:0] adc1_p, adc1_n,
    input wire data_clock_p, data_clock_n,
    input wire frame_clock_p, frame_clock_n,
    output wire adc_ref_clock_p, adc_ref_clock_n,   //this one is the reference for the sampling
    //spi interface
    input wire adc_sdo,
    output wire adc_sdi,
    output wire adc_cs_n,
    output wire adc_sck,

    //ADC data
    output wire adc_clock,
    output wire [15:0] adc0_data, adc1_data,
    output wire adc_data_valid,
    output wire idelay_rdy
);

//we dont use the spi 
assign adc_sdi = 1;
assign adc_cs_n = 1;
assign adc_sck = 1;

generate
    //only if the fpga geneartes the sampling clock
    if(OUTPUT_CLOCK)begin
    output_clock output_clock_inst (
        .clk(clk),
        .adc_ref_clk_p(adc_ref_clock_p),
        .adc_ref_clk_n(adc_ref_clock_n)
    );
    end
endgenerate


//create clokcs 
wire data_clk_bufio, data_clk_div;
wire iserdes2_bitslip;          //this one is generated by the clock alignment and used in the data_phy also
wire [2:0] bitslip_count;
reg sync_rst=0; //this one is set a little bit ahead
wire frame_valid;


clock_alignment #(
    .IOSTANDARD(IOSTANDARD),
    .BUFR_DIVIDE(BUFR_DIVIDE_CLOCK)
) clock_alignment_inst (
    .data_clock_p(data_clock_p),
    .data_clock_n(data_clock_n),
    .frame_clock_p(frame_clock_p),
    .frame_clock_n(frame_clock_n),
    .async_rst(async_rst),
    .sync_rst(sync_rst),
    .data_clk_bufio(data_clk_bufio),
    .data_clk_div(data_clk_div),
    .frame_valid(frame_valid),
    .iserdes2_bitslip(iserdes2_bitslip),
    .bitslip_count(bitslip_count)
);

//logic reset
//serdes rst should be held at least two cycles
reg [7:0] serdes_rst_cnt=16;
always@(posedge data_clk_div or posedge async_rst)begin
    if(async_rst)begin
        sync_rst = 1;
        serdes_rst_cnt <= 16;
    end
    else begin
        if(serdes_rst_cnt >0)begin
            serdes_rst_cnt <= serdes_rst_cnt-1;
            sync_rst <= 1;
        end
        else 
            sync_rst <= 0;
    end
end

//idealyctrl reset, should be held for T_IDELAYCTRL_RPW (60ns) after configuration 
//with the a 200mhz reference should be held 12 cycles minimum
reg idelay_rst;
reg [7:0] idelay_rst_cnt=16;
always@(posedge idelay_ref)begin
    if(async_rst)begin
        idelay_rst_cnt <= 16;
        idelay_rst<=1;
    end
    else begin
        if(idelay_rst_cnt>0)begin
            idelay_rst_cnt <= idelay_rst_cnt-1;
            idelay_rst <= 1;
        end
        else
            idelay_rst <= 0;
    end
end

//instantiate idelayctrl
IDELAYCTRL idelay_adc (
	.RST    (idelay_rst),
	.REFCLK (idelay_ref),
	.RDY    (idelay_rdy)
);

//data phy

data_phy #(
    .ARCH(ARCHITECTURE)
) data_phy_adc [1:0] ( 
    .sync_rst(sync_rst), 
    .adc_data_p({adc0_p, adc1_p}), 
    .adc_data_n({adc0_n, adc1_n}),
    .data_clk_bufio(data_clk_bufio),
    .data_clk_div(data_clk_div),
    .bitslip(iserdes2_bitslip),
    .adc_data({adc0_data, adc1_data})
);


assign adc_clock = data_clk_div;
assign adc_data_valid = frame_valid;

endmodule
