`default_nettype none

module complex_add #(
    parameter DIN_WIDTH = 32,
    parameter DIN_POINT = 
    pa


)
