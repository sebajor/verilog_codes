`default_nettype none
`include "agc.v"


module agc_tb #(
    parameter DIN_WIDTH = 8,    //its ufix8_7
    parameter DELAY_LINE = 32,
    parameter REFRESH_CYCLES = 1024,
    parameter GAIN_WIDTH = 12,   //its ufix12_10
    parameter [GAIN_WIDTH-1:0] GAIN_LOW_LIM = 12'd12    //the gain couldnt be less than this
) (
    input wire clk,
    input wire rst,

    input wire signed [DIN_WIDTH-1:0] din,
    input wire din_valid,
    
    input wire [2*DIN_WIDTH-1:0] ref_pow,    //ufix16_14    reference power
    input wire [2*DIN_WIDTH-1:0] error_coef, //ufix16_14    coef to adjust the error
                                             //before adding it to the gain

    output wire [DIN_WIDTH-1:0] dout,
    output wire dout_valid
);


agc #(
    .DIN_WIDTH(DIN_WIDTH),
    .DELAY_LINE(DELAY_LINE),
    .REFRESH_CYCLES(REFRESH_CYCLES),
    .GAIN_WIDTH(GAIN_WIDTH),
    .GAIN_LOW_LIM(GAIN_LOW_LIM)
) agc_inst (
    .clk(clk),
    .rst(rst),
    .din(din),
    .din_valid(din_valid),
    .ref_pow(ref_pow),    
    .error_coef(error_coef),
    .dout(dout),
    .dout_valid(dout_valid)
);

initial begin
    $dumpfile("traces.vcd");
    $dumpvars();
end


endmodule
