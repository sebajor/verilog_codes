`default_nettype none
`include "includes.v"


module r22sdf_fft16 #(
    parameter DIN_WIDTH = 16,
    parameter DIN_POINT = 14,
    parameter TWIDD_WIDTH = 16,
    parameter 


)
