`default_nettype none

module acc_ctrl #(
    parameter 


)
