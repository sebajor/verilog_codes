`default_nettype none
`include "rtl/sync_simple_dual_ram.v"

module unsign_vacc #(
    parameter DIN_WIDTH = 32,
    parameter VECTOR_LEN = 64,
    parameter DOUT_WIDTH = 64
) (
    input wire clk,
    input wire new_acc,     //new accumulation, set it previous the first sample of the frame
    
    input wire [DIN_WIDTH-1:0] din,
    input wire din_valid,

    output wire [DOUT_WIDTH-1:0] dout,
    output wire dout_valid
);

reg [$clog2(VECTOR_LEN)-1:0] w_addr=0, r_addr=1;
reg [$clog2(VECTOR_LEN):0] acc_count=0;
reg [2*DIN_WIDTH-1:0] din_r=0;
reg [2:0] din_valid_r=0;
reg add_zero=0;
reg [1:0] add_zero_r=0;

always@(posedge clk)begin
    din_valid_r <= {din_valid_r[1:0], din_valid};
    din_r <= {din_r[DIN_WIDTH-1:0], din};
    add_zero_r <= {add_zero_r[0], add_zero};
    if(new_acc)
        add_zero <= 1'b1;
    else if(add_zero & (acc_count == (VECTOR_LEN-1)) & din_valid)
        add_zero <= 1'b0;
end


//pointers logic
always@(posedge clk)begin
    if(din_valid)begin
        r_addr <= r_addr+1;
        if(add_zero)begin
            if(acc_count == (VECTOR_LEN-1))
                acc_count <=0;
            else
                acc_count <= acc_count+1;
        end
        else
            acc_count <=0;
    end
    if(din_valid_r[2])
        w_addr<= w_addr+1;
end

wire [DOUT_WIDTH-1:0] bram_out;
reg [DOUT_WIDTH-1:0] acc=0;

sync_simple_dual_ram #(
    .RAM_WIDTH(DOUT_WIDTH),
    .RAM_DEPTH(VECTOR_LEN),
    .RAM_PERFORMANCE("HIGH_PERFORMANCE")
) ram_inst  (
    .clka(clk),
    .addra(w_addr),
    .dina(acc),
    .wea(din_valid_r[2]),   //check!!!
    .addrb(r_addr),
    .enb(1'b1),
    .rstb(1'b0), 
    .regceb(1'b1),
    .doutb(bram_out)         // RAM output data
);

reg [2*DOUT_WIDTH-1:0] bram_out_r=0;
always@(posedge clk)begin
    if(din_valid_r[0])
        bram_out_r <= {bram_out_r[DOUT_WIDTH-1:0], bram_out};
end


wire [DOUT_WIDTH-1:0] actual_acc = bram_out_r[2*DOUT_WIDTH-1:DOUT_WIDTH];

reg dout_valid_r=0;
wire [DIN_WIDTH-1:0] din_delay = din_r[DIN_WIDTH+:DIN_WIDTH];

always@(posedge clk)begin
    if(din_valid_r[1])begin
        if(add_zero_r[1])begin
            acc <= din_delay;
            dout_valid_r <=1;
            //acc_count <= acc_count+1;
        end
        else begin
            acc <= actual_acc+din_delay;
            dout_valid_r <=0;
            //acc_count <=0;
        end
    end
    else 
        dout_valid_r <=0;
end


assign dout = actual_acc;//bram_out;
assign dout_valid = dout_valid_r;




endmodule
