`default_nettype none

module dvi #(


)
